-------------------------------------------------------------------------------
-- lmb_bram_elaborate.vhd
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

entity lmb_bram_elaborate is
  generic (
    C_MEMSIZE : integer;
    C_PORT_DWIDTH : integer;
    C_PORT_AWIDTH : integer;
    C_NUM_WE : integer;
    C_FAMILY : string
    );
  port (
    BRAM_Rst_A : in std_logic;
    BRAM_Clk_A : in std_logic;
    BRAM_EN_A : in std_logic;
    BRAM_WEN_A : in std_logic_vector(0 to C_NUM_WE-1);
    BRAM_Addr_A : in std_logic_vector(0 to C_PORT_AWIDTH-1);
    BRAM_Din_A : out std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Dout_A : in std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Rst_B : in std_logic;
    BRAM_Clk_B : in std_logic;
    BRAM_EN_B : in std_logic;
    BRAM_WEN_B : in std_logic_vector(0 to C_NUM_WE-1);
    BRAM_Addr_B : in std_logic_vector(0 to C_PORT_AWIDTH-1);
    BRAM_Din_B : out std_logic_vector(0 to C_PORT_DWIDTH-1);
    BRAM_Dout_B : in std_logic_vector(0 to C_PORT_DWIDTH-1)
  );

  attribute keep_hierarchy : STRING;
  attribute keep_hierarchy of lmb_bram_elaborate : entity is "yes";

end lmb_bram_elaborate;

architecture STRUCTURE of lmb_bram_elaborate is

  component RAMB36 is
    generic (
      WRITE_MODE_A : string;
      WRITE_MODE_B : string;
      READ_WIDTH_A : integer;
      READ_WIDTH_B : integer;
      WRITE_WIDTH_A : integer;
      WRITE_WIDTH_B : integer;
      RAM_EXTENSION_A : string;
      RAM_EXTENSION_B : string
    );
    port (
      ADDRA : in std_logic_vector(15 downto 0);
      CASCADEINLATA : in std_logic;
      CASCADEINREGA : in std_logic;
      CASCADEOUTLATA : out std_logic;
      CASCADEOUTREGA : out std_logic;
      CLKA : in std_logic;
      DIA : in std_logic_vector(31 downto 0);
      DIPA : in std_logic_vector(3 downto 0);
      DOA : out std_logic_vector(31 downto 0);
      DOPA : out std_logic_vector(3 downto 0);
      ENA : in std_logic;
      REGCEA : in std_logic;
      SSRA : in std_logic;
      WEA : in std_logic_vector(3 downto 0);
      ADDRB : in std_logic_vector(15 downto 0);
      CASCADEINLATB : in std_logic;
      CASCADEINREGB : in std_logic;
      CASCADEOUTLATB : out std_logic;
      CASCADEOUTREGB : out std_logic;
      CLKB : in std_logic;
      DIB : in std_logic_vector(31 downto 0);
      DIPB : in std_logic_vector(3 downto 0);
      DOB : out std_logic_vector(31 downto 0);
      DOPB : out std_logic_vector(3 downto 0);
      ENB : in std_logic;
      REGCEB : in std_logic;
      SSRB : in std_logic;
      WEB : in std_logic_vector(3 downto 0)
    );
  end component;

  -- Internal signals

  signal net_gnd0 : std_logic;
  signal net_gnd4 : std_logic_vector(3 downto 0);
  signal pgassign1 : std_logic_vector(0 to 0);
  signal pgassign2 : std_logic_vector(0 to 30);
  signal pgassign3 : std_logic_vector(15 downto 0);
  signal pgassign4 : std_logic_vector(31 downto 0);
  signal pgassign5 : std_logic_vector(31 downto 0);
  signal pgassign6 : std_logic_vector(3 downto 0);
  signal pgassign7 : std_logic_vector(15 downto 0);
  signal pgassign8 : std_logic_vector(31 downto 0);
  signal pgassign9 : std_logic_vector(31 downto 0);
  signal pgassign10 : std_logic_vector(3 downto 0);
  signal pgassign11 : std_logic_vector(15 downto 0);
  signal pgassign12 : std_logic_vector(31 downto 0);
  signal pgassign13 : std_logic_vector(31 downto 0);
  signal pgassign14 : std_logic_vector(3 downto 0);
  signal pgassign15 : std_logic_vector(15 downto 0);
  signal pgassign16 : std_logic_vector(31 downto 0);
  signal pgassign17 : std_logic_vector(31 downto 0);
  signal pgassign18 : std_logic_vector(3 downto 0);
  signal pgassign19 : std_logic_vector(15 downto 0);
  signal pgassign20 : std_logic_vector(31 downto 0);
  signal pgassign21 : std_logic_vector(31 downto 0);
  signal pgassign22 : std_logic_vector(3 downto 0);
  signal pgassign23 : std_logic_vector(15 downto 0);
  signal pgassign24 : std_logic_vector(31 downto 0);
  signal pgassign25 : std_logic_vector(31 downto 0);
  signal pgassign26 : std_logic_vector(3 downto 0);
  signal pgassign27 : std_logic_vector(15 downto 0);
  signal pgassign28 : std_logic_vector(31 downto 0);
  signal pgassign29 : std_logic_vector(31 downto 0);
  signal pgassign30 : std_logic_vector(3 downto 0);
  signal pgassign31 : std_logic_vector(15 downto 0);
  signal pgassign32 : std_logic_vector(31 downto 0);
  signal pgassign33 : std_logic_vector(31 downto 0);
  signal pgassign34 : std_logic_vector(3 downto 0);
  signal pgassign35 : std_logic_vector(15 downto 0);
  signal pgassign36 : std_logic_vector(31 downto 0);
  signal pgassign37 : std_logic_vector(31 downto 0);
  signal pgassign38 : std_logic_vector(3 downto 0);
  signal pgassign39 : std_logic_vector(15 downto 0);
  signal pgassign40 : std_logic_vector(31 downto 0);
  signal pgassign41 : std_logic_vector(31 downto 0);
  signal pgassign42 : std_logic_vector(3 downto 0);
  signal pgassign43 : std_logic_vector(15 downto 0);
  signal pgassign44 : std_logic_vector(31 downto 0);
  signal pgassign45 : std_logic_vector(31 downto 0);
  signal pgassign46 : std_logic_vector(3 downto 0);
  signal pgassign47 : std_logic_vector(15 downto 0);
  signal pgassign48 : std_logic_vector(31 downto 0);
  signal pgassign49 : std_logic_vector(31 downto 0);
  signal pgassign50 : std_logic_vector(3 downto 0);
  signal pgassign51 : std_logic_vector(15 downto 0);
  signal pgassign52 : std_logic_vector(31 downto 0);
  signal pgassign53 : std_logic_vector(31 downto 0);
  signal pgassign54 : std_logic_vector(3 downto 0);
  signal pgassign55 : std_logic_vector(15 downto 0);
  signal pgassign56 : std_logic_vector(31 downto 0);
  signal pgassign57 : std_logic_vector(31 downto 0);
  signal pgassign58 : std_logic_vector(3 downto 0);
  signal pgassign59 : std_logic_vector(15 downto 0);
  signal pgassign60 : std_logic_vector(31 downto 0);
  signal pgassign61 : std_logic_vector(31 downto 0);
  signal pgassign62 : std_logic_vector(3 downto 0);
  signal pgassign63 : std_logic_vector(15 downto 0);
  signal pgassign64 : std_logic_vector(31 downto 0);
  signal pgassign65 : std_logic_vector(31 downto 0);
  signal pgassign66 : std_logic_vector(3 downto 0);
  signal pgassign67 : std_logic_vector(15 downto 0);
  signal pgassign68 : std_logic_vector(31 downto 0);
  signal pgassign69 : std_logic_vector(31 downto 0);
  signal pgassign70 : std_logic_vector(3 downto 0);
  signal pgassign71 : std_logic_vector(15 downto 0);
  signal pgassign72 : std_logic_vector(31 downto 0);
  signal pgassign73 : std_logic_vector(31 downto 0);
  signal pgassign74 : std_logic_vector(3 downto 0);
  signal pgassign75 : std_logic_vector(15 downto 0);
  signal pgassign76 : std_logic_vector(31 downto 0);
  signal pgassign77 : std_logic_vector(31 downto 0);
  signal pgassign78 : std_logic_vector(3 downto 0);
  signal pgassign79 : std_logic_vector(15 downto 0);
  signal pgassign80 : std_logic_vector(31 downto 0);
  signal pgassign81 : std_logic_vector(31 downto 0);
  signal pgassign82 : std_logic_vector(3 downto 0);
  signal pgassign83 : std_logic_vector(15 downto 0);
  signal pgassign84 : std_logic_vector(31 downto 0);
  signal pgassign85 : std_logic_vector(31 downto 0);
  signal pgassign86 : std_logic_vector(3 downto 0);
  signal pgassign87 : std_logic_vector(15 downto 0);
  signal pgassign88 : std_logic_vector(31 downto 0);
  signal pgassign89 : std_logic_vector(31 downto 0);
  signal pgassign90 : std_logic_vector(3 downto 0);
  signal pgassign91 : std_logic_vector(15 downto 0);
  signal pgassign92 : std_logic_vector(31 downto 0);
  signal pgassign93 : std_logic_vector(31 downto 0);
  signal pgassign94 : std_logic_vector(3 downto 0);
  signal pgassign95 : std_logic_vector(15 downto 0);
  signal pgassign96 : std_logic_vector(31 downto 0);
  signal pgassign97 : std_logic_vector(31 downto 0);
  signal pgassign98 : std_logic_vector(3 downto 0);
  signal pgassign99 : std_logic_vector(15 downto 0);
  signal pgassign100 : std_logic_vector(31 downto 0);
  signal pgassign101 : std_logic_vector(31 downto 0);
  signal pgassign102 : std_logic_vector(3 downto 0);
  signal pgassign103 : std_logic_vector(15 downto 0);
  signal pgassign104 : std_logic_vector(31 downto 0);
  signal pgassign105 : std_logic_vector(31 downto 0);
  signal pgassign106 : std_logic_vector(3 downto 0);
  signal pgassign107 : std_logic_vector(15 downto 0);
  signal pgassign108 : std_logic_vector(31 downto 0);
  signal pgassign109 : std_logic_vector(31 downto 0);
  signal pgassign110 : std_logic_vector(3 downto 0);
  signal pgassign111 : std_logic_vector(15 downto 0);
  signal pgassign112 : std_logic_vector(31 downto 0);
  signal pgassign113 : std_logic_vector(31 downto 0);
  signal pgassign114 : std_logic_vector(3 downto 0);
  signal pgassign115 : std_logic_vector(15 downto 0);
  signal pgassign116 : std_logic_vector(31 downto 0);
  signal pgassign117 : std_logic_vector(31 downto 0);
  signal pgassign118 : std_logic_vector(3 downto 0);
  signal pgassign119 : std_logic_vector(15 downto 0);
  signal pgassign120 : std_logic_vector(31 downto 0);
  signal pgassign121 : std_logic_vector(31 downto 0);
  signal pgassign122 : std_logic_vector(3 downto 0);
  signal pgassign123 : std_logic_vector(15 downto 0);
  signal pgassign124 : std_logic_vector(31 downto 0);
  signal pgassign125 : std_logic_vector(31 downto 0);
  signal pgassign126 : std_logic_vector(3 downto 0);
  signal pgassign127 : std_logic_vector(15 downto 0);
  signal pgassign128 : std_logic_vector(31 downto 0);
  signal pgassign129 : std_logic_vector(31 downto 0);
  signal pgassign130 : std_logic_vector(3 downto 0);
  signal pgassign131 : std_logic_vector(15 downto 0);
  signal pgassign132 : std_logic_vector(31 downto 0);
  signal pgassign133 : std_logic_vector(31 downto 0);
  signal pgassign134 : std_logic_vector(3 downto 0);
  signal pgassign135 : std_logic_vector(15 downto 0);
  signal pgassign136 : std_logic_vector(31 downto 0);
  signal pgassign137 : std_logic_vector(31 downto 0);
  signal pgassign138 : std_logic_vector(3 downto 0);
  signal pgassign139 : std_logic_vector(15 downto 0);
  signal pgassign140 : std_logic_vector(31 downto 0);
  signal pgassign141 : std_logic_vector(31 downto 0);
  signal pgassign142 : std_logic_vector(3 downto 0);
  signal pgassign143 : std_logic_vector(15 downto 0);
  signal pgassign144 : std_logic_vector(31 downto 0);
  signal pgassign145 : std_logic_vector(31 downto 0);
  signal pgassign146 : std_logic_vector(3 downto 0);
  signal pgassign147 : std_logic_vector(15 downto 0);
  signal pgassign148 : std_logic_vector(31 downto 0);
  signal pgassign149 : std_logic_vector(31 downto 0);
  signal pgassign150 : std_logic_vector(3 downto 0);
  signal pgassign151 : std_logic_vector(15 downto 0);
  signal pgassign152 : std_logic_vector(31 downto 0);
  signal pgassign153 : std_logic_vector(31 downto 0);
  signal pgassign154 : std_logic_vector(3 downto 0);
  signal pgassign155 : std_logic_vector(15 downto 0);
  signal pgassign156 : std_logic_vector(31 downto 0);
  signal pgassign157 : std_logic_vector(31 downto 0);
  signal pgassign158 : std_logic_vector(3 downto 0);
  signal pgassign159 : std_logic_vector(15 downto 0);
  signal pgassign160 : std_logic_vector(31 downto 0);
  signal pgassign161 : std_logic_vector(31 downto 0);
  signal pgassign162 : std_logic_vector(3 downto 0);
  signal pgassign163 : std_logic_vector(15 downto 0);
  signal pgassign164 : std_logic_vector(31 downto 0);
  signal pgassign165 : std_logic_vector(31 downto 0);
  signal pgassign166 : std_logic_vector(3 downto 0);
  signal pgassign167 : std_logic_vector(15 downto 0);
  signal pgassign168 : std_logic_vector(31 downto 0);
  signal pgassign169 : std_logic_vector(31 downto 0);
  signal pgassign170 : std_logic_vector(3 downto 0);
  signal pgassign171 : std_logic_vector(15 downto 0);
  signal pgassign172 : std_logic_vector(31 downto 0);
  signal pgassign173 : std_logic_vector(31 downto 0);
  signal pgassign174 : std_logic_vector(3 downto 0);
  signal pgassign175 : std_logic_vector(15 downto 0);
  signal pgassign176 : std_logic_vector(31 downto 0);
  signal pgassign177 : std_logic_vector(31 downto 0);
  signal pgassign178 : std_logic_vector(3 downto 0);
  signal pgassign179 : std_logic_vector(15 downto 0);
  signal pgassign180 : std_logic_vector(31 downto 0);
  signal pgassign181 : std_logic_vector(31 downto 0);
  signal pgassign182 : std_logic_vector(3 downto 0);
  signal pgassign183 : std_logic_vector(15 downto 0);
  signal pgassign184 : std_logic_vector(31 downto 0);
  signal pgassign185 : std_logic_vector(31 downto 0);
  signal pgassign186 : std_logic_vector(3 downto 0);
  signal pgassign187 : std_logic_vector(15 downto 0);
  signal pgassign188 : std_logic_vector(31 downto 0);
  signal pgassign189 : std_logic_vector(31 downto 0);
  signal pgassign190 : std_logic_vector(3 downto 0);
  signal pgassign191 : std_logic_vector(15 downto 0);
  signal pgassign192 : std_logic_vector(31 downto 0);
  signal pgassign193 : std_logic_vector(31 downto 0);
  signal pgassign194 : std_logic_vector(3 downto 0);
  signal pgassign195 : std_logic_vector(15 downto 0);
  signal pgassign196 : std_logic_vector(31 downto 0);
  signal pgassign197 : std_logic_vector(31 downto 0);
  signal pgassign198 : std_logic_vector(3 downto 0);
  signal pgassign199 : std_logic_vector(15 downto 0);
  signal pgassign200 : std_logic_vector(31 downto 0);
  signal pgassign201 : std_logic_vector(31 downto 0);
  signal pgassign202 : std_logic_vector(3 downto 0);
  signal pgassign203 : std_logic_vector(15 downto 0);
  signal pgassign204 : std_logic_vector(31 downto 0);
  signal pgassign205 : std_logic_vector(31 downto 0);
  signal pgassign206 : std_logic_vector(3 downto 0);
  signal pgassign207 : std_logic_vector(15 downto 0);
  signal pgassign208 : std_logic_vector(31 downto 0);
  signal pgassign209 : std_logic_vector(31 downto 0);
  signal pgassign210 : std_logic_vector(3 downto 0);
  signal pgassign211 : std_logic_vector(15 downto 0);
  signal pgassign212 : std_logic_vector(31 downto 0);
  signal pgassign213 : std_logic_vector(31 downto 0);
  signal pgassign214 : std_logic_vector(3 downto 0);
  signal pgassign215 : std_logic_vector(15 downto 0);
  signal pgassign216 : std_logic_vector(31 downto 0);
  signal pgassign217 : std_logic_vector(31 downto 0);
  signal pgassign218 : std_logic_vector(3 downto 0);
  signal pgassign219 : std_logic_vector(15 downto 0);
  signal pgassign220 : std_logic_vector(31 downto 0);
  signal pgassign221 : std_logic_vector(31 downto 0);
  signal pgassign222 : std_logic_vector(3 downto 0);
  signal pgassign223 : std_logic_vector(15 downto 0);
  signal pgassign224 : std_logic_vector(31 downto 0);
  signal pgassign225 : std_logic_vector(31 downto 0);
  signal pgassign226 : std_logic_vector(3 downto 0);
  signal pgassign227 : std_logic_vector(15 downto 0);
  signal pgassign228 : std_logic_vector(31 downto 0);
  signal pgassign229 : std_logic_vector(31 downto 0);
  signal pgassign230 : std_logic_vector(3 downto 0);
  signal pgassign231 : std_logic_vector(15 downto 0);
  signal pgassign232 : std_logic_vector(31 downto 0);
  signal pgassign233 : std_logic_vector(31 downto 0);
  signal pgassign234 : std_logic_vector(3 downto 0);
  signal pgassign235 : std_logic_vector(15 downto 0);
  signal pgassign236 : std_logic_vector(31 downto 0);
  signal pgassign237 : std_logic_vector(31 downto 0);
  signal pgassign238 : std_logic_vector(3 downto 0);
  signal pgassign239 : std_logic_vector(15 downto 0);
  signal pgassign240 : std_logic_vector(31 downto 0);
  signal pgassign241 : std_logic_vector(31 downto 0);
  signal pgassign242 : std_logic_vector(3 downto 0);
  signal pgassign243 : std_logic_vector(15 downto 0);
  signal pgassign244 : std_logic_vector(31 downto 0);
  signal pgassign245 : std_logic_vector(31 downto 0);
  signal pgassign246 : std_logic_vector(3 downto 0);
  signal pgassign247 : std_logic_vector(15 downto 0);
  signal pgassign248 : std_logic_vector(31 downto 0);
  signal pgassign249 : std_logic_vector(31 downto 0);
  signal pgassign250 : std_logic_vector(3 downto 0);
  signal pgassign251 : std_logic_vector(15 downto 0);
  signal pgassign252 : std_logic_vector(31 downto 0);
  signal pgassign253 : std_logic_vector(31 downto 0);
  signal pgassign254 : std_logic_vector(3 downto 0);
  signal pgassign255 : std_logic_vector(15 downto 0);
  signal pgassign256 : std_logic_vector(31 downto 0);
  signal pgassign257 : std_logic_vector(31 downto 0);
  signal pgassign258 : std_logic_vector(3 downto 0);

begin

  -- Internal assignments

  pgassign1(0 to 0) <= B"1";
  pgassign2(0 to 30) <= B"0000000000000000000000000000000";
  pgassign3(15 downto 15) <= B"1";
  pgassign3(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign4(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign4(0 downto 0) <= BRAM_Dout_A(0 to 0);
  BRAM_Din_A(0 to 0) <= pgassign5(0 downto 0);
  pgassign6(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign6(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign6(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign6(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign7(15 downto 15) <= B"1";
  pgassign7(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign8(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign8(0 downto 0) <= BRAM_Dout_B(0 to 0);
  BRAM_Din_B(0 to 0) <= pgassign9(0 downto 0);
  pgassign10(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign10(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign10(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign10(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign11(15 downto 15) <= B"1";
  pgassign11(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign12(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign12(0 downto 0) <= BRAM_Dout_A(1 to 1);
  BRAM_Din_A(1 to 1) <= pgassign13(0 downto 0);
  pgassign14(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign14(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign14(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign14(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign15(15 downto 15) <= B"1";
  pgassign15(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign16(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign16(0 downto 0) <= BRAM_Dout_B(1 to 1);
  BRAM_Din_B(1 to 1) <= pgassign17(0 downto 0);
  pgassign18(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign18(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign18(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign18(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign19(15 downto 15) <= B"1";
  pgassign19(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign20(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign20(0 downto 0) <= BRAM_Dout_A(2 to 2);
  BRAM_Din_A(2 to 2) <= pgassign21(0 downto 0);
  pgassign22(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign22(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign22(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign22(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign23(15 downto 15) <= B"1";
  pgassign23(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign24(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign24(0 downto 0) <= BRAM_Dout_B(2 to 2);
  BRAM_Din_B(2 to 2) <= pgassign25(0 downto 0);
  pgassign26(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign26(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign26(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign26(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign27(15 downto 15) <= B"1";
  pgassign27(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign28(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign28(0 downto 0) <= BRAM_Dout_A(3 to 3);
  BRAM_Din_A(3 to 3) <= pgassign29(0 downto 0);
  pgassign30(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign30(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign30(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign30(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign31(15 downto 15) <= B"1";
  pgassign31(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign32(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign32(0 downto 0) <= BRAM_Dout_B(3 to 3);
  BRAM_Din_B(3 to 3) <= pgassign33(0 downto 0);
  pgassign34(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign34(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign34(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign34(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign35(15 downto 15) <= B"1";
  pgassign35(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign36(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign36(0 downto 0) <= BRAM_Dout_A(4 to 4);
  BRAM_Din_A(4 to 4) <= pgassign37(0 downto 0);
  pgassign38(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign38(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign38(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign38(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign39(15 downto 15) <= B"1";
  pgassign39(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign40(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign40(0 downto 0) <= BRAM_Dout_B(4 to 4);
  BRAM_Din_B(4 to 4) <= pgassign41(0 downto 0);
  pgassign42(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign42(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign42(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign42(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign43(15 downto 15) <= B"1";
  pgassign43(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign44(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign44(0 downto 0) <= BRAM_Dout_A(5 to 5);
  BRAM_Din_A(5 to 5) <= pgassign45(0 downto 0);
  pgassign46(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign46(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign46(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign46(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign47(15 downto 15) <= B"1";
  pgassign47(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign48(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign48(0 downto 0) <= BRAM_Dout_B(5 to 5);
  BRAM_Din_B(5 to 5) <= pgassign49(0 downto 0);
  pgassign50(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign50(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign50(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign50(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign51(15 downto 15) <= B"1";
  pgassign51(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign52(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign52(0 downto 0) <= BRAM_Dout_A(6 to 6);
  BRAM_Din_A(6 to 6) <= pgassign53(0 downto 0);
  pgassign54(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign54(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign54(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign54(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign55(15 downto 15) <= B"1";
  pgassign55(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign56(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign56(0 downto 0) <= BRAM_Dout_B(6 to 6);
  BRAM_Din_B(6 to 6) <= pgassign57(0 downto 0);
  pgassign58(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign58(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign58(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign58(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign59(15 downto 15) <= B"1";
  pgassign59(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign60(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign60(0 downto 0) <= BRAM_Dout_A(7 to 7);
  BRAM_Din_A(7 to 7) <= pgassign61(0 downto 0);
  pgassign62(3 downto 3) <= BRAM_WEN_A(0 to 0);
  pgassign62(2 downto 2) <= BRAM_WEN_A(0 to 0);
  pgassign62(1 downto 1) <= BRAM_WEN_A(0 to 0);
  pgassign62(0 downto 0) <= BRAM_WEN_A(0 to 0);
  pgassign63(15 downto 15) <= B"1";
  pgassign63(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign64(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign64(0 downto 0) <= BRAM_Dout_B(7 to 7);
  BRAM_Din_B(7 to 7) <= pgassign65(0 downto 0);
  pgassign66(3 downto 3) <= BRAM_WEN_B(0 to 0);
  pgassign66(2 downto 2) <= BRAM_WEN_B(0 to 0);
  pgassign66(1 downto 1) <= BRAM_WEN_B(0 to 0);
  pgassign66(0 downto 0) <= BRAM_WEN_B(0 to 0);
  pgassign67(15 downto 15) <= B"1";
  pgassign67(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign68(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign68(0 downto 0) <= BRAM_Dout_A(8 to 8);
  BRAM_Din_A(8 to 8) <= pgassign69(0 downto 0);
  pgassign70(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign70(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign70(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign70(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign71(15 downto 15) <= B"1";
  pgassign71(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign72(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign72(0 downto 0) <= BRAM_Dout_B(8 to 8);
  BRAM_Din_B(8 to 8) <= pgassign73(0 downto 0);
  pgassign74(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign74(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign74(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign74(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign75(15 downto 15) <= B"1";
  pgassign75(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign76(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign76(0 downto 0) <= BRAM_Dout_A(9 to 9);
  BRAM_Din_A(9 to 9) <= pgassign77(0 downto 0);
  pgassign78(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign78(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign78(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign78(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign79(15 downto 15) <= B"1";
  pgassign79(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign80(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign80(0 downto 0) <= BRAM_Dout_B(9 to 9);
  BRAM_Din_B(9 to 9) <= pgassign81(0 downto 0);
  pgassign82(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign82(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign82(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign82(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign83(15 downto 15) <= B"1";
  pgassign83(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign84(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign84(0 downto 0) <= BRAM_Dout_A(10 to 10);
  BRAM_Din_A(10 to 10) <= pgassign85(0 downto 0);
  pgassign86(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign86(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign86(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign86(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign87(15 downto 15) <= B"1";
  pgassign87(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign88(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign88(0 downto 0) <= BRAM_Dout_B(10 to 10);
  BRAM_Din_B(10 to 10) <= pgassign89(0 downto 0);
  pgassign90(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign90(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign90(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign90(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign91(15 downto 15) <= B"1";
  pgassign91(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign92(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign92(0 downto 0) <= BRAM_Dout_A(11 to 11);
  BRAM_Din_A(11 to 11) <= pgassign93(0 downto 0);
  pgassign94(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign94(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign94(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign94(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign95(15 downto 15) <= B"1";
  pgassign95(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign96(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign96(0 downto 0) <= BRAM_Dout_B(11 to 11);
  BRAM_Din_B(11 to 11) <= pgassign97(0 downto 0);
  pgassign98(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign98(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign98(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign98(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign99(15 downto 15) <= B"1";
  pgassign99(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign100(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign100(0 downto 0) <= BRAM_Dout_A(12 to 12);
  BRAM_Din_A(12 to 12) <= pgassign101(0 downto 0);
  pgassign102(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign102(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign102(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign102(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign103(15 downto 15) <= B"1";
  pgassign103(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign104(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign104(0 downto 0) <= BRAM_Dout_B(12 to 12);
  BRAM_Din_B(12 to 12) <= pgassign105(0 downto 0);
  pgassign106(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign106(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign106(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign106(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign107(15 downto 15) <= B"1";
  pgassign107(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign108(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign108(0 downto 0) <= BRAM_Dout_A(13 to 13);
  BRAM_Din_A(13 to 13) <= pgassign109(0 downto 0);
  pgassign110(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign110(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign110(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign110(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign111(15 downto 15) <= B"1";
  pgassign111(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign112(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign112(0 downto 0) <= BRAM_Dout_B(13 to 13);
  BRAM_Din_B(13 to 13) <= pgassign113(0 downto 0);
  pgassign114(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign114(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign114(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign114(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign115(15 downto 15) <= B"1";
  pgassign115(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign116(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign116(0 downto 0) <= BRAM_Dout_A(14 to 14);
  BRAM_Din_A(14 to 14) <= pgassign117(0 downto 0);
  pgassign118(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign118(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign118(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign118(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign119(15 downto 15) <= B"1";
  pgassign119(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign120(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign120(0 downto 0) <= BRAM_Dout_B(14 to 14);
  BRAM_Din_B(14 to 14) <= pgassign121(0 downto 0);
  pgassign122(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign122(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign122(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign122(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign123(15 downto 15) <= B"1";
  pgassign123(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign124(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign124(0 downto 0) <= BRAM_Dout_A(15 to 15);
  BRAM_Din_A(15 to 15) <= pgassign125(0 downto 0);
  pgassign126(3 downto 3) <= BRAM_WEN_A(1 to 1);
  pgassign126(2 downto 2) <= BRAM_WEN_A(1 to 1);
  pgassign126(1 downto 1) <= BRAM_WEN_A(1 to 1);
  pgassign126(0 downto 0) <= BRAM_WEN_A(1 to 1);
  pgassign127(15 downto 15) <= B"1";
  pgassign127(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign128(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign128(0 downto 0) <= BRAM_Dout_B(15 to 15);
  BRAM_Din_B(15 to 15) <= pgassign129(0 downto 0);
  pgassign130(3 downto 3) <= BRAM_WEN_B(1 to 1);
  pgassign130(2 downto 2) <= BRAM_WEN_B(1 to 1);
  pgassign130(1 downto 1) <= BRAM_WEN_B(1 to 1);
  pgassign130(0 downto 0) <= BRAM_WEN_B(1 to 1);
  pgassign131(15 downto 15) <= B"1";
  pgassign131(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign132(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign132(0 downto 0) <= BRAM_Dout_A(16 to 16);
  BRAM_Din_A(16 to 16) <= pgassign133(0 downto 0);
  pgassign134(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign134(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign134(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign134(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign135(15 downto 15) <= B"1";
  pgassign135(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign136(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign136(0 downto 0) <= BRAM_Dout_B(16 to 16);
  BRAM_Din_B(16 to 16) <= pgassign137(0 downto 0);
  pgassign138(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign138(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign138(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign138(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign139(15 downto 15) <= B"1";
  pgassign139(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign140(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign140(0 downto 0) <= BRAM_Dout_A(17 to 17);
  BRAM_Din_A(17 to 17) <= pgassign141(0 downto 0);
  pgassign142(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign142(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign142(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign142(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign143(15 downto 15) <= B"1";
  pgassign143(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign144(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign144(0 downto 0) <= BRAM_Dout_B(17 to 17);
  BRAM_Din_B(17 to 17) <= pgassign145(0 downto 0);
  pgassign146(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign146(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign146(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign146(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign147(15 downto 15) <= B"1";
  pgassign147(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign148(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign148(0 downto 0) <= BRAM_Dout_A(18 to 18);
  BRAM_Din_A(18 to 18) <= pgassign149(0 downto 0);
  pgassign150(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign150(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign150(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign150(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign151(15 downto 15) <= B"1";
  pgassign151(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign152(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign152(0 downto 0) <= BRAM_Dout_B(18 to 18);
  BRAM_Din_B(18 to 18) <= pgassign153(0 downto 0);
  pgassign154(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign154(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign154(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign154(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign155(15 downto 15) <= B"1";
  pgassign155(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign156(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign156(0 downto 0) <= BRAM_Dout_A(19 to 19);
  BRAM_Din_A(19 to 19) <= pgassign157(0 downto 0);
  pgassign158(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign158(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign158(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign158(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign159(15 downto 15) <= B"1";
  pgassign159(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign160(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign160(0 downto 0) <= BRAM_Dout_B(19 to 19);
  BRAM_Din_B(19 to 19) <= pgassign161(0 downto 0);
  pgassign162(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign162(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign162(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign162(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign163(15 downto 15) <= B"1";
  pgassign163(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign164(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign164(0 downto 0) <= BRAM_Dout_A(20 to 20);
  BRAM_Din_A(20 to 20) <= pgassign165(0 downto 0);
  pgassign166(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign166(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign166(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign166(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign167(15 downto 15) <= B"1";
  pgassign167(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign168(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign168(0 downto 0) <= BRAM_Dout_B(20 to 20);
  BRAM_Din_B(20 to 20) <= pgassign169(0 downto 0);
  pgassign170(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign170(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign170(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign170(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign171(15 downto 15) <= B"1";
  pgassign171(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign172(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign172(0 downto 0) <= BRAM_Dout_A(21 to 21);
  BRAM_Din_A(21 to 21) <= pgassign173(0 downto 0);
  pgassign174(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign174(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign174(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign174(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign175(15 downto 15) <= B"1";
  pgassign175(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign176(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign176(0 downto 0) <= BRAM_Dout_B(21 to 21);
  BRAM_Din_B(21 to 21) <= pgassign177(0 downto 0);
  pgassign178(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign178(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign178(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign178(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign179(15 downto 15) <= B"1";
  pgassign179(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign180(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign180(0 downto 0) <= BRAM_Dout_A(22 to 22);
  BRAM_Din_A(22 to 22) <= pgassign181(0 downto 0);
  pgassign182(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign182(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign182(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign182(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign183(15 downto 15) <= B"1";
  pgassign183(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign184(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign184(0 downto 0) <= BRAM_Dout_B(22 to 22);
  BRAM_Din_B(22 to 22) <= pgassign185(0 downto 0);
  pgassign186(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign186(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign186(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign186(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign187(15 downto 15) <= B"1";
  pgassign187(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign188(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign188(0 downto 0) <= BRAM_Dout_A(23 to 23);
  BRAM_Din_A(23 to 23) <= pgassign189(0 downto 0);
  pgassign190(3 downto 3) <= BRAM_WEN_A(2 to 2);
  pgassign190(2 downto 2) <= BRAM_WEN_A(2 to 2);
  pgassign190(1 downto 1) <= BRAM_WEN_A(2 to 2);
  pgassign190(0 downto 0) <= BRAM_WEN_A(2 to 2);
  pgassign191(15 downto 15) <= B"1";
  pgassign191(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign192(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign192(0 downto 0) <= BRAM_Dout_B(23 to 23);
  BRAM_Din_B(23 to 23) <= pgassign193(0 downto 0);
  pgassign194(3 downto 3) <= BRAM_WEN_B(2 to 2);
  pgassign194(2 downto 2) <= BRAM_WEN_B(2 to 2);
  pgassign194(1 downto 1) <= BRAM_WEN_B(2 to 2);
  pgassign194(0 downto 0) <= BRAM_WEN_B(2 to 2);
  pgassign195(15 downto 15) <= B"1";
  pgassign195(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign196(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign196(0 downto 0) <= BRAM_Dout_A(24 to 24);
  BRAM_Din_A(24 to 24) <= pgassign197(0 downto 0);
  pgassign198(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign198(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign198(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign198(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign199(15 downto 15) <= B"1";
  pgassign199(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign200(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign200(0 downto 0) <= BRAM_Dout_B(24 to 24);
  BRAM_Din_B(24 to 24) <= pgassign201(0 downto 0);
  pgassign202(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign202(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign202(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign202(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign203(15 downto 15) <= B"1";
  pgassign203(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign204(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign204(0 downto 0) <= BRAM_Dout_A(25 to 25);
  BRAM_Din_A(25 to 25) <= pgassign205(0 downto 0);
  pgassign206(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign206(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign206(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign206(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign207(15 downto 15) <= B"1";
  pgassign207(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign208(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign208(0 downto 0) <= BRAM_Dout_B(25 to 25);
  BRAM_Din_B(25 to 25) <= pgassign209(0 downto 0);
  pgassign210(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign210(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign210(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign210(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign211(15 downto 15) <= B"1";
  pgassign211(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign212(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign212(0 downto 0) <= BRAM_Dout_A(26 to 26);
  BRAM_Din_A(26 to 26) <= pgassign213(0 downto 0);
  pgassign214(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign214(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign214(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign214(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign215(15 downto 15) <= B"1";
  pgassign215(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign216(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign216(0 downto 0) <= BRAM_Dout_B(26 to 26);
  BRAM_Din_B(26 to 26) <= pgassign217(0 downto 0);
  pgassign218(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign218(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign218(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign218(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign219(15 downto 15) <= B"1";
  pgassign219(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign220(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign220(0 downto 0) <= BRAM_Dout_A(27 to 27);
  BRAM_Din_A(27 to 27) <= pgassign221(0 downto 0);
  pgassign222(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign222(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign222(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign222(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign223(15 downto 15) <= B"1";
  pgassign223(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign224(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign224(0 downto 0) <= BRAM_Dout_B(27 to 27);
  BRAM_Din_B(27 to 27) <= pgassign225(0 downto 0);
  pgassign226(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign226(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign226(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign226(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign227(15 downto 15) <= B"1";
  pgassign227(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign228(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign228(0 downto 0) <= BRAM_Dout_A(28 to 28);
  BRAM_Din_A(28 to 28) <= pgassign229(0 downto 0);
  pgassign230(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign230(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign230(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign230(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign231(15 downto 15) <= B"1";
  pgassign231(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign232(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign232(0 downto 0) <= BRAM_Dout_B(28 to 28);
  BRAM_Din_B(28 to 28) <= pgassign233(0 downto 0);
  pgassign234(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign234(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign234(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign234(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign235(15 downto 15) <= B"1";
  pgassign235(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign236(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign236(0 downto 0) <= BRAM_Dout_A(29 to 29);
  BRAM_Din_A(29 to 29) <= pgassign237(0 downto 0);
  pgassign238(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign238(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign238(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign238(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign239(15 downto 15) <= B"1";
  pgassign239(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign240(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign240(0 downto 0) <= BRAM_Dout_B(29 to 29);
  BRAM_Din_B(29 to 29) <= pgassign241(0 downto 0);
  pgassign242(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign242(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign242(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign242(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign243(15 downto 15) <= B"1";
  pgassign243(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign244(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign244(0 downto 0) <= BRAM_Dout_A(30 to 30);
  BRAM_Din_A(30 to 30) <= pgassign245(0 downto 0);
  pgassign246(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign246(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign246(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign246(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign247(15 downto 15) <= B"1";
  pgassign247(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign248(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign248(0 downto 0) <= BRAM_Dout_B(30 to 30);
  BRAM_Din_B(30 to 30) <= pgassign249(0 downto 0);
  pgassign250(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign250(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign250(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign250(0 downto 0) <= BRAM_WEN_B(3 to 3);
  pgassign251(15 downto 15) <= B"1";
  pgassign251(14 downto 0) <= BRAM_Addr_A(15 to 29);
  pgassign252(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign252(0 downto 0) <= BRAM_Dout_A(31 to 31);
  BRAM_Din_A(31 to 31) <= pgassign253(0 downto 0);
  pgassign254(3 downto 3) <= BRAM_WEN_A(3 to 3);
  pgassign254(2 downto 2) <= BRAM_WEN_A(3 to 3);
  pgassign254(1 downto 1) <= BRAM_WEN_A(3 to 3);
  pgassign254(0 downto 0) <= BRAM_WEN_A(3 to 3);
  pgassign255(15 downto 15) <= B"1";
  pgassign255(14 downto 0) <= BRAM_Addr_B(15 to 29);
  pgassign256(31 downto 1) <= B"0000000000000000000000000000000";
  pgassign256(0 downto 0) <= BRAM_Dout_B(31 to 31);
  BRAM_Din_B(31 to 31) <= pgassign257(0 downto 0);
  pgassign258(3 downto 3) <= BRAM_WEN_B(3 to 3);
  pgassign258(2 downto 2) <= BRAM_WEN_B(3 to 3);
  pgassign258(1 downto 1) <= BRAM_WEN_B(3 to 3);
  pgassign258(0 downto 0) <= BRAM_WEN_B(3 to 3);
  net_gnd0 <= '0';
  net_gnd4(3 downto 0) <= B"0000";

  ramb36_0 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign3,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign4,
      DIPA => net_gnd4,
      DOA => pgassign5,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign6,
      ADDRB => pgassign7,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign8,
      DIPB => net_gnd4,
      DOB => pgassign9,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign10
    );

  ramb36_1 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign11,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign12,
      DIPA => net_gnd4,
      DOA => pgassign13,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign14,
      ADDRB => pgassign15,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign16,
      DIPB => net_gnd4,
      DOB => pgassign17,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign18
    );

  ramb36_2 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign19,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign20,
      DIPA => net_gnd4,
      DOA => pgassign21,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign22,
      ADDRB => pgassign23,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign24,
      DIPB => net_gnd4,
      DOB => pgassign25,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign26
    );

  ramb36_3 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign27,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign28,
      DIPA => net_gnd4,
      DOA => pgassign29,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign30,
      ADDRB => pgassign31,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign32,
      DIPB => net_gnd4,
      DOB => pgassign33,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign34
    );

  ramb36_4 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign35,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign36,
      DIPA => net_gnd4,
      DOA => pgassign37,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign38,
      ADDRB => pgassign39,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign40,
      DIPB => net_gnd4,
      DOB => pgassign41,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign42
    );

  ramb36_5 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign43,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign44,
      DIPA => net_gnd4,
      DOA => pgassign45,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign46,
      ADDRB => pgassign47,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign48,
      DIPB => net_gnd4,
      DOB => pgassign49,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign50
    );

  ramb36_6 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign51,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign52,
      DIPA => net_gnd4,
      DOA => pgassign53,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign54,
      ADDRB => pgassign55,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign56,
      DIPB => net_gnd4,
      DOB => pgassign57,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign58
    );

  ramb36_7 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign59,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign60,
      DIPA => net_gnd4,
      DOA => pgassign61,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign62,
      ADDRB => pgassign63,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign64,
      DIPB => net_gnd4,
      DOB => pgassign65,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign66
    );

  ramb36_8 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign67,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign68,
      DIPA => net_gnd4,
      DOA => pgassign69,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign70,
      ADDRB => pgassign71,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign72,
      DIPB => net_gnd4,
      DOB => pgassign73,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign74
    );

  ramb36_9 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign75,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign76,
      DIPA => net_gnd4,
      DOA => pgassign77,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign78,
      ADDRB => pgassign79,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign80,
      DIPB => net_gnd4,
      DOB => pgassign81,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign82
    );

  ramb36_10 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign83,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign84,
      DIPA => net_gnd4,
      DOA => pgassign85,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign86,
      ADDRB => pgassign87,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign88,
      DIPB => net_gnd4,
      DOB => pgassign89,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign90
    );

  ramb36_11 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign91,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign92,
      DIPA => net_gnd4,
      DOA => pgassign93,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign94,
      ADDRB => pgassign95,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign96,
      DIPB => net_gnd4,
      DOB => pgassign97,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign98
    );

  ramb36_12 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign99,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign100,
      DIPA => net_gnd4,
      DOA => pgassign101,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign102,
      ADDRB => pgassign103,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign104,
      DIPB => net_gnd4,
      DOB => pgassign105,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign106
    );

  ramb36_13 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign107,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign108,
      DIPA => net_gnd4,
      DOA => pgassign109,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign110,
      ADDRB => pgassign111,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign112,
      DIPB => net_gnd4,
      DOB => pgassign113,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign114
    );

  ramb36_14 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign115,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign116,
      DIPA => net_gnd4,
      DOA => pgassign117,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign118,
      ADDRB => pgassign119,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign120,
      DIPB => net_gnd4,
      DOB => pgassign121,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign122
    );

  ramb36_15 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign123,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign124,
      DIPA => net_gnd4,
      DOA => pgassign125,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign126,
      ADDRB => pgassign127,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign128,
      DIPB => net_gnd4,
      DOB => pgassign129,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign130
    );

  ramb36_16 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign131,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign132,
      DIPA => net_gnd4,
      DOA => pgassign133,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign134,
      ADDRB => pgassign135,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign136,
      DIPB => net_gnd4,
      DOB => pgassign137,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign138
    );

  ramb36_17 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign139,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign140,
      DIPA => net_gnd4,
      DOA => pgassign141,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign142,
      ADDRB => pgassign143,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign144,
      DIPB => net_gnd4,
      DOB => pgassign145,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign146
    );

  ramb36_18 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign147,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign148,
      DIPA => net_gnd4,
      DOA => pgassign149,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign150,
      ADDRB => pgassign151,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign152,
      DIPB => net_gnd4,
      DOB => pgassign153,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign154
    );

  ramb36_19 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign155,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign156,
      DIPA => net_gnd4,
      DOA => pgassign157,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign158,
      ADDRB => pgassign159,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign160,
      DIPB => net_gnd4,
      DOB => pgassign161,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign162
    );

  ramb36_20 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign163,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign164,
      DIPA => net_gnd4,
      DOA => pgassign165,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign166,
      ADDRB => pgassign167,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign168,
      DIPB => net_gnd4,
      DOB => pgassign169,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign170
    );

  ramb36_21 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign171,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign172,
      DIPA => net_gnd4,
      DOA => pgassign173,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign174,
      ADDRB => pgassign175,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign176,
      DIPB => net_gnd4,
      DOB => pgassign177,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign178
    );

  ramb36_22 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign179,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign180,
      DIPA => net_gnd4,
      DOA => pgassign181,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign182,
      ADDRB => pgassign183,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign184,
      DIPB => net_gnd4,
      DOB => pgassign185,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign186
    );

  ramb36_23 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign187,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign188,
      DIPA => net_gnd4,
      DOA => pgassign189,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign190,
      ADDRB => pgassign191,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign192,
      DIPB => net_gnd4,
      DOB => pgassign193,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign194
    );

  ramb36_24 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign195,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign196,
      DIPA => net_gnd4,
      DOA => pgassign197,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign198,
      ADDRB => pgassign199,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign200,
      DIPB => net_gnd4,
      DOB => pgassign201,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign202
    );

  ramb36_25 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign203,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign204,
      DIPA => net_gnd4,
      DOA => pgassign205,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign206,
      ADDRB => pgassign207,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign208,
      DIPB => net_gnd4,
      DOB => pgassign209,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign210
    );

  ramb36_26 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign211,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign212,
      DIPA => net_gnd4,
      DOA => pgassign213,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign214,
      ADDRB => pgassign215,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign216,
      DIPB => net_gnd4,
      DOB => pgassign217,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign218
    );

  ramb36_27 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign219,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign220,
      DIPA => net_gnd4,
      DOA => pgassign221,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign222,
      ADDRB => pgassign223,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign224,
      DIPB => net_gnd4,
      DOB => pgassign225,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign226
    );

  ramb36_28 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign227,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign228,
      DIPA => net_gnd4,
      DOA => pgassign229,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign230,
      ADDRB => pgassign231,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign232,
      DIPB => net_gnd4,
      DOB => pgassign233,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign234
    );

  ramb36_29 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign235,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign236,
      DIPA => net_gnd4,
      DOA => pgassign237,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign238,
      ADDRB => pgassign239,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign240,
      DIPB => net_gnd4,
      DOB => pgassign241,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign242
    );

  ramb36_30 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign243,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign244,
      DIPA => net_gnd4,
      DOA => pgassign245,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign246,
      ADDRB => pgassign247,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign248,
      DIPB => net_gnd4,
      DOB => pgassign249,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign250
    );

  ramb36_31 : RAMB36
    generic map (
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      READ_WIDTH_A => 1,
      READ_WIDTH_B => 1,
      WRITE_WIDTH_A => 1,
      WRITE_WIDTH_B => 1,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE"
    )
    port map (
      ADDRA => pgassign251,
      CASCADEINLATA => net_gnd0,
      CASCADEINREGA => net_gnd0,
      CASCADEOUTLATA => open,
      CASCADEOUTREGA => open,
      CLKA => BRAM_Clk_A,
      DIA => pgassign252,
      DIPA => net_gnd4,
      DOA => pgassign253,
      DOPA => open,
      ENA => BRAM_EN_A,
      REGCEA => net_gnd0,
      SSRA => BRAM_Rst_A,
      WEA => pgassign254,
      ADDRB => pgassign255,
      CASCADEINLATB => net_gnd0,
      CASCADEINREGB => net_gnd0,
      CASCADEOUTLATB => open,
      CASCADEOUTREGB => open,
      CLKB => BRAM_Clk_B,
      DIB => pgassign256,
      DIPB => net_gnd4,
      DOB => pgassign257,
      DOPB => open,
      ENB => BRAM_EN_B,
      REGCEB => net_gnd0,
      SSRB => BRAM_Rst_B,
      WEB => pgassign258
    );

end architecture STRUCTURE;

